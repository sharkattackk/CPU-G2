`timescale 1ns / 1ns
// XOR module

module XOR(m, x, y);
    input x, y;
    outputm;

    assign m = x ^ y;  
endmodule