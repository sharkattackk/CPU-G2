module rotate_right(
output [31:0] R,
input [31:0] A, B
);

	wire [4:0] M;
	assign M = A % 32;
	assign R = (M == 31) ? {B[30:0], B[31:31]} :

												(M == 30) ? {B[29:0], B[31:30]} :
												(M == 29) ? {B[28:0], B[31:29]} :
												(M == 28) ? {B[27:0], B[31:28]} :
												(M == 27) ? {B[26:0], B[31:27]} :
												(M == 26) ? {B[25:0], B[31:26]} :
												(M == 25) ? {B[24:0], B[31:25]} :
												(M == 24) ? {B[23:0], B[31:24]} :
												(M == 23) ? {B[22:0], B[31:23]} :
												(M == 22) ? {B[21:0], B[31:22]} :
												(M == 21) ? {B[20:0], B[31:21]} :
												(M == 20) ? {B[19:0], B[31:20]} :
												(M == 19) ? {B[18:0], B[31:19]} :
												(M == 18) ? {B[17:0], B[31:18]} :
												(M == 17) ? {B[16:0], B[31:17]} :
												(M == 16) ? {B[15:0], B[31:16]} :
												(M == 15) ? {B[14:0], B[31:15]} :
												(M == 14) ? {B[13:0], B[31:14]} :
												(M == 13) ? {B[12:0], B[31:13]} :
												(M == 12) ? {B[11:0], B[31:12]} :
												(M == 11) ? {B[10:0], B[31:11]} :
												(M == 10) ? {B[9:0], B[31:10]} :
												(M == 9) ? {B[8:0], B[31:9]} :
												(M == 8) ? {B[7:0], B[31:8]} :
												(M == 7) ? {B[6:0], B[31:7]} :
												(M == 6) ? {B[5:0], B[31:6]} :
												(M == 5) ? {B[4:0], B[31:5]} :
												(M == 4) ? {B[3:0], B[31:4]} :
												(M == 3) ? {B[2:0], B[31:3]} :
												(M == 2) ? {B[1:0], B[31:2]} :
												(M == 1) ? {B[0:0], B[31:1]} :
												 B[31:0];
endmodule