`timescale 1ns / 1ns
// OR module

module OR(cOut, x, y);
    input [31:0] x, y;
    output [31:0] m;

    m = x | y;  
endmodule