`timescale 1ns / 1ns
// Booths Algorithm Module
module MUL(M, Q, P);
    input [31:0] M, Q;
    output reg [63:0] P;

    
